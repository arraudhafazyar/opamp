magic
tech sky130A
magscale 1 2
timestamp 1729166590
<< nwell >>
rect -176 -1526 1008 1439
<< nsubdiff >>
rect -140 1369 -80 1403
rect 896 1369 956 1403
rect -140 1347 -106 1369
rect 922 1347 956 1369
rect -140 -1456 -106 -1434
rect 922 -1456 956 -1434
rect -140 -1490 -80 -1456
rect 896 -1490 956 -1456
<< nsubdiffcont >>
rect -80 1369 896 1403
rect -140 -1434 -106 1347
rect 922 -1434 956 1347
rect -80 -1490 896 -1456
<< poly >>
rect -56 1319 36 1335
rect -56 1285 -40 1319
rect -6 1285 36 1319
rect -56 1269 36 1285
rect 6 1264 36 1269
rect 610 1319 702 1335
rect 610 1285 652 1319
rect 686 1285 702 1319
rect 610 1269 702 1285
rect 610 1260 640 1269
rect 94 641 295 741
rect -56 625 36 641
rect -56 591 -40 625
rect -6 591 36 625
rect -56 575 36 591
rect 6 570 36 575
rect 610 625 702 641
rect 610 591 652 625
rect 686 591 702 625
rect 610 575 702 591
rect 610 570 640 575
rect 94 45 294 47
rect 352 45 553 48
rect 93 -53 553 45
rect 93 -55 551 -53
rect 6 -581 36 -575
rect -56 -597 36 -581
rect -56 -631 -40 -597
rect -6 -631 36 -597
rect -56 -647 36 -631
rect 610 -581 640 -576
rect 610 -597 702 -581
rect 610 -631 652 -597
rect 686 -631 702 -597
rect 352 -745 552 -646
rect 610 -647 702 -631
rect 6 -1273 36 -1267
rect -56 -1289 36 -1273
rect -56 -1323 -40 -1289
rect -6 -1323 36 -1289
rect -56 -1339 36 -1323
rect 610 -1273 640 -1267
rect 610 -1289 702 -1273
rect 610 -1323 652 -1289
rect 686 -1323 702 -1289
rect 610 -1339 702 -1323
<< polycont >>
rect -40 1285 -6 1319
rect 652 1285 686 1319
rect -40 591 -6 625
rect 652 591 686 625
rect -40 -631 -6 -597
rect 652 -631 686 -597
rect -40 -1323 -6 -1289
rect 652 -1323 686 -1289
<< locali >>
rect -140 1369 -80 1403
rect 896 1369 956 1403
rect -140 1347 -106 1369
rect 922 1347 956 1369
rect -56 1285 -40 1319
rect -6 1285 10 1319
rect 636 1285 652 1319
rect 686 1285 702 1319
rect -40 1221 -6 1285
rect 652 1201 686 1285
rect -56 591 -40 625
rect -6 591 10 625
rect 636 591 652 625
rect 686 591 702 625
rect -40 512 -5 591
rect 652 508 686 591
rect -40 -597 -6 -510
rect 652 -597 686 -518
rect -56 -631 -40 -597
rect -6 -631 10 -597
rect 636 -631 652 -597
rect 686 -631 702 -597
rect -40 -1289 -6 -1221
rect 652 -1289 687 -1209
rect -56 -1323 -40 -1289
rect -6 -1323 10 -1289
rect 636 -1323 652 -1289
rect 686 -1323 702 -1289
rect -140 -1456 -106 -1434
rect 922 -1456 956 -1434
rect -140 -1490 -80 -1456
rect 896 -1490 956 -1456
<< viali >>
rect 652 1369 686 1403
rect -40 1285 -6 1319
rect 652 1285 686 1319
rect -40 591 -6 625
rect 652 591 686 625
rect -40 -631 -6 -597
rect 652 -631 686 -597
rect -40 -1323 -6 -1289
rect 652 -1323 686 -1289
rect -40 -1490 -6 -1456
<< metal1 >>
rect 640 1403 698 1409
rect 640 1369 652 1403
rect 686 1369 698 1403
rect 640 1359 698 1369
rect -52 1319 6 1325
rect -52 1285 -40 1319
rect -6 1285 6 1319
rect -52 1279 6 1285
rect 640 1319 699 1359
rect 640 1285 652 1319
rect 686 1285 699 1319
rect 640 1283 699 1285
rect 640 1279 698 1283
rect -50 1228 6 1279
rect -59 849 -49 1228
rect 3 1226 13 1228
rect 3 850 73 1226
rect 3 849 13 850
rect 300 797 346 1238
rect 646 1226 695 1279
rect 571 1194 695 1226
rect 571 850 677 1194
rect 558 797 604 838
rect 300 751 383 797
rect 523 751 604 797
rect -52 625 6 631
rect -52 591 -40 625
rect -6 591 6 625
rect -52 585 6 591
rect -49 534 0 585
rect 28 531 38 535
rect -34 155 38 531
rect 91 155 101 535
rect 44 -109 198 -63
rect 44 -163 90 -109
rect -34 -164 90 -163
rect -34 -514 72 -164
rect -52 -539 72 -514
rect -52 -591 4 -539
rect -52 -597 6 -591
rect -52 -631 -40 -597
rect -6 -631 6 -597
rect -52 -637 6 -631
rect 300 -759 346 751
rect 640 625 698 631
rect 640 591 652 625
rect 686 591 698 625
rect 640 585 698 591
rect 644 570 695 585
rect 644 532 692 570
rect 573 506 692 532
rect 573 156 679 506
rect 564 97 598 156
rect 504 63 598 97
rect 546 -537 556 -162
rect 608 -518 679 -162
rect 608 -537 695 -518
rect 573 -538 695 -537
rect 646 -591 695 -538
rect 640 -597 698 -591
rect 640 -631 652 -597
rect 686 -631 698 -597
rect 640 -637 698 -631
rect 42 -796 130 -760
rect 42 -855 78 -796
rect 252 -797 346 -759
rect -32 -886 78 -855
rect -32 -1214 74 -886
rect -49 -1231 74 -1214
rect -49 -1283 0 -1231
rect 300 -1242 346 -797
rect 633 -855 643 -853
rect 578 -1231 643 -855
rect 633 -1233 643 -1231
rect 695 -1233 705 -853
rect 646 -1283 695 -1233
rect -52 -1289 6 -1283
rect -52 -1323 -40 -1289
rect -6 -1323 6 -1289
rect -52 -1456 6 -1323
rect 640 -1289 698 -1283
rect 640 -1323 652 -1289
rect 686 -1323 698 -1289
rect 640 -1329 698 -1323
rect -52 -1490 -40 -1456
rect -6 -1490 6 -1456
rect -52 -1496 6 -1490
<< via1 >>
rect -49 849 3 1228
rect 38 155 91 535
rect 556 -537 608 -162
rect 643 -1233 695 -853
<< metal2 >>
rect -49 1229 3 1238
rect -50 1228 3 1229
rect -50 850 -49 1228
rect -49 735 3 849
rect 641 735 697 742
rect -62 675 -53 735
rect 7 675 16 735
rect 639 733 699 735
rect 639 677 641 733
rect 697 677 699 733
rect -50 -648 -2 675
rect 38 535 91 545
rect 38 145 91 155
rect 40 106 90 145
rect 40 37 89 106
rect 40 -12 607 37
rect 558 -152 607 -12
rect 556 -162 608 -152
rect 556 -547 608 -537
rect -54 -657 2 -648
rect 639 -655 699 677
rect -54 -722 2 -713
rect 630 -715 639 -655
rect 699 -715 708 -655
rect 639 -853 699 -715
rect 639 -892 643 -853
rect 695 -892 699 -853
rect 643 -1243 695 -1233
<< via2 >>
rect -53 675 7 735
rect 641 677 697 733
rect -54 -713 2 -657
rect 639 -715 699 -655
<< metal3 >>
rect -58 735 12 740
rect 636 735 702 738
rect -58 675 -53 735
rect 7 733 702 735
rect 7 677 641 733
rect 697 677 702 733
rect 7 675 702 677
rect -58 670 12 675
rect 636 672 702 675
rect -59 -655 7 -652
rect 634 -655 704 -650
rect -59 -657 639 -655
rect -59 -713 -54 -657
rect 2 -713 639 -657
rect -59 -715 639 -713
rect 699 -715 704 -655
rect -59 -718 7 -715
rect 634 -720 704 -715
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729135466
transform 1 0 625 0 1 -1042
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729135466
transform 1 0 21 0 1 -1042
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729135466
transform 1 0 625 0 1 344
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729135466
transform 1 0 21 0 1 -350
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729135466
transform 1 0 625 0 1 -350
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729135466
transform 1 0 21 0 1 344
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729135466
transform 1 0 625 0 1 1038
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729135466
transform 1 0 21 0 1 1038
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729138823
transform 1 0 323 0 1 1038
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729138823
transform 1 0 323 0 1 344
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729138823
transform 1 0 323 0 1 -350
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729138823
transform 1 0 323 0 1 -1042
box -323 -300 323 300
<< labels >>
flabel metal1 667 1348 667 1348 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal2 62 77 62 77 0 FreeSans 160 0 0 0 D1
port 1 nsew
flabel metal1 582 108 585 109 0 FreeSans 160 0 0 0 D2
port 2 nsew
flabel metal2 673 61 673 61 0 FreeSans 160 0 0 0 D5
port 3 nsew
<< end >>
