magic
tech sky130A
magscale 1 2
timestamp 1729428391
<< dnwell >>
rect -10 2016 2104 4050
<< nwell >>
rect -63 1963 2157 4103
<< viali >>
rect 939 2895 1094 2931
rect 1249 2903 1285 3027
rect 1662 488 1760 524
rect 1998 336 2096 388
<< metal1 >>
rect 1243 3037 1291 3039
rect 925 3027 1291 3037
rect 925 2931 1249 3027
rect 925 2895 939 2931
rect 1094 2903 1249 2931
rect 1285 2903 1291 3027
rect 1094 2895 1291 2903
rect 1420 2896 1421 2958
rect 925 2891 1291 2895
rect 925 2888 1284 2891
rect 1317 1627 1323 1634
rect 740 1589 1323 1627
rect 1317 1582 1323 1589
rect 1375 1582 1381 1634
rect 719 1509 729 1561
rect 783 1509 1260 1561
rect 1208 1281 1260 1509
rect 1208 1229 1656 1281
rect 1651 530 1661 534
rect 1650 482 1661 530
rect 1759 530 1769 534
rect 1759 524 1772 530
rect 1760 488 1772 524
rect 1759 482 1772 488
rect 1986 388 2108 394
rect 1986 336 1998 388
rect 2096 336 2108 388
rect 1986 330 2108 336
rect 2606 -85 2658 -79
rect 2401 -135 2606 -89
rect 2606 -143 2658 -137
<< via1 >>
rect 1323 1582 1375 1634
rect 729 1509 783 1561
rect 1661 524 1759 534
rect 1661 488 1662 524
rect 1662 488 1759 524
rect 1661 482 1759 488
rect 1998 336 2096 388
rect 2606 -137 2658 -85
<< metal2 >>
rect 1714 2566 1766 2594
rect 1886 2219 2525 2261
rect 1330 1831 1549 1869
rect 1330 1640 1368 1831
rect 1511 1763 1549 1831
rect 1323 1634 1375 1640
rect 1323 1576 1375 1582
rect 729 1561 783 1571
rect 729 1499 783 1509
rect 1661 534 1759 544
rect 1640 482 1661 523
rect 1759 482 2161 523
rect 1640 388 2161 482
rect 2483 470 2525 2219
rect 2602 2177 2662 2186
rect 2602 2108 2662 2117
rect 1640 337 1998 388
rect 2096 337 2161 388
rect 2320 428 2525 470
rect 1998 326 2096 336
rect 2320 231 2362 428
rect 2609 -85 2655 2108
rect 2600 -137 2606 -85
rect 2658 -137 2664 -85
<< via2 >>
rect 2602 2117 2662 2177
<< metal3 >>
rect 1305 2579 1693 2641
rect 1305 2262 1367 2579
rect 800 2200 1367 2262
rect 2597 2177 2667 2182
rect 1794 2117 2602 2177
rect 2662 2117 2667 2177
rect 2597 2112 2667 2117
rect 1865 1283 1927 1310
rect 1755 1109 1822 1129
use differential  differential_0
timestamp 1729408613
transform 1 0 1437 0 1 3495
box -223 -1479 668 554
use nmoscs2  nmoscs2_0
timestamp 1729241942
transform 1 0 1435 0 1 -456
box -176 -165 1106 851
use nmoscs  nmoscs_0
timestamp 1729408613
transform 1 0 1497 0 1 1227
box -229 -744 908 711
use pmoscs  pmoscs_0
timestamp 1729166590
transform 1 0 176 0 1 1526
box -176 -1526 1008 1439
<< labels >>
flabel metal2 1913 443 1913 443 0 FreeSans 1600 0 0 0 gnd
port 5 nsew
flabel metal2 2418 2238 2418 2238 0 FreeSans 320 0 0 0 out
port 7 nsew
flabel metal2 1734 2578 1734 2578 0 FreeSans 320 0 0 0 vpin
port 8 nsew
flabel nwell 1580 3486 1580 3486 0 FreeSans 320 0 0 0 vin
port 9 nsew
flabel metal3 1895 1296 1895 1296 0 FreeSans 320 0 0 0 rs
port 10 nsew
flabel metal1 1125 2966 1125 2966 0 FreeSans 320 0 0 0 vdd
port 12 nsew
<< end >>
