magic
tech sky130A
magscale 1 2
timestamp 1729408613
<< nwell >>
rect -223 -1479 668 554
<< nsubdiff >>
rect -187 484 -127 518
rect 572 484 632 518
rect -187 462 -153 484
rect 598 462 632 484
rect -187 -1409 -153 -1383
rect 598 -1409 632 -1383
rect -187 -1443 -127 -1409
rect 572 -1443 632 -1409
<< nsubdiffcont >>
rect -127 484 572 518
rect -187 -1383 -153 462
rect 598 -1383 632 462
rect -127 -1443 572 -1409
<< poly >>
rect 6 69 36 75
rect -56 53 36 69
rect -56 19 -40 53
rect -6 19 36 53
rect -56 3 36 19
rect 410 69 440 88
rect 410 53 501 69
rect 410 19 451 53
rect 485 19 501 53
rect 410 3 501 19
rect -56 -108 36 -92
rect -56 -142 -40 -108
rect -6 -142 36 -108
rect -56 -158 36 -142
rect 6 -175 36 -158
rect 410 -108 502 -92
rect 410 -142 452 -108
rect 486 -142 502 -108
rect 410 -158 502 -142
rect 410 -175 440 -158
rect 6 -759 36 -746
rect 415 -753 440 -752
rect -56 -775 36 -759
rect -56 -809 -40 -775
rect -6 -809 36 -775
rect -56 -825 36 -809
rect 410 -760 440 -753
rect 410 -776 501 -760
rect 410 -810 451 -776
rect 485 -810 501 -776
rect 410 -826 501 -810
rect -55 -945 37 -929
rect -55 -979 -39 -945
rect -5 -979 37 -945
rect -55 -995 37 -979
rect 7 -1000 37 -995
rect 411 -945 503 -929
rect 411 -979 453 -945
rect 487 -979 503 -945
rect 411 -995 503 -979
rect 411 -1000 441 -995
<< polycont >>
rect -40 19 -6 53
rect 451 19 485 53
rect -40 -142 -6 -108
rect 452 -142 486 -108
rect -40 -809 -6 -775
rect 451 -810 485 -776
rect -39 -979 -5 -945
rect 453 -979 487 -945
<< locali >>
rect -187 484 -127 518
rect 572 484 632 518
rect -187 462 -153 484
rect 598 462 632 484
rect -40 53 -6 129
rect 451 53 485 136
rect -56 19 -40 53
rect -6 19 10 53
rect 435 19 451 53
rect 485 19 501 53
rect 452 -108 486 -107
rect -56 -142 -40 -108
rect -6 -142 10 -108
rect 436 -142 452 -108
rect 486 -142 502 -108
rect -40 -229 -6 -142
rect 452 -231 486 -142
rect -40 -775 -6 -697
rect -56 -809 -40 -775
rect -6 -809 10 -775
rect 451 -776 486 -699
rect -40 -810 -6 -809
rect 435 -810 451 -776
rect 485 -810 501 -776
rect -55 -979 -39 -945
rect -5 -979 11 -945
rect 437 -979 453 -945
rect 487 -979 503 -945
rect -39 -1067 -5 -979
rect 453 -1063 487 -979
rect -187 -1409 -153 -1383
rect 598 -1409 632 -1383
rect -187 -1443 -127 -1409
rect 572 -1443 632 -1409
<< viali >>
rect 24 518 179 523
rect 24 484 179 518
rect 24 483 179 484
rect -40 19 -6 53
rect 451 19 485 53
rect -40 -142 -6 -108
rect 452 -142 486 -108
rect -40 -809 -6 -775
rect 451 -810 485 -776
rect -39 -979 -5 -945
rect 453 -979 487 -945
<< metal1 >>
rect 12 523 191 529
rect 12 483 24 523
rect 179 483 191 523
rect 12 477 191 483
rect -37 129 39 300
rect -46 101 39 129
rect 91 101 101 300
rect -46 59 -2 101
rect 185 100 195 301
rect 251 100 261 301
rect 368 100 442 300
rect 494 100 504 300
rect -52 53 6 59
rect 121 53 166 59
rect -52 19 -40 53
rect -6 19 6 53
rect 110 19 178 53
rect -52 13 6 19
rect 121 -31 166 19
rect 266 10 276 62
rect 328 10 338 62
rect 445 59 489 100
rect 439 53 497 59
rect 439 19 451 53
rect 485 19 497 53
rect 439 13 497 19
rect 121 -76 325 -31
rect -52 -108 6 -102
rect -52 -142 -40 -108
rect -6 -142 6 -108
rect -52 -148 6 -142
rect -46 -200 0 -148
rect 108 -162 118 -110
rect 170 -162 180 -110
rect 280 -159 325 -76
rect 440 -108 498 -102
rect 440 -142 452 -108
rect 486 -142 498 -108
rect 440 -148 498 -142
rect 447 -199 490 -148
rect -59 -401 -49 -200
rect 3 -400 75 -200
rect 185 -400 195 -200
rect 251 -400 261 -200
rect 346 -400 356 -199
rect 408 -237 490 -199
rect 408 -400 481 -237
rect 3 -401 13 -400
rect -59 -728 -49 -527
rect 3 -728 79 -527
rect 367 -528 482 -527
rect 185 -728 195 -528
rect 251 -728 261 -528
rect 345 -728 355 -528
rect 407 -699 482 -528
rect 407 -728 491 -699
rect -47 -769 0 -728
rect -52 -775 6 -769
rect -52 -809 -40 -775
rect -6 -809 6 -775
rect -52 -815 6 -809
rect 107 -818 117 -766
rect 169 -818 179 -766
rect 283 -857 328 -769
rect 445 -770 491 -728
rect 439 -776 497 -770
rect 439 -810 451 -776
rect 485 -810 497 -776
rect 439 -816 497 -810
rect 124 -902 328 -857
rect -51 -945 7 -939
rect -51 -979 -39 -945
rect -5 -979 7 -945
rect -51 -985 7 -979
rect 124 -985 169 -902
rect 267 -985 277 -933
rect 329 -985 339 -933
rect 441 -945 499 -939
rect 441 -979 453 -945
rect 487 -979 499 -945
rect 441 -985 499 -979
rect -43 -1026 -1 -985
rect 448 -1024 492 -985
rect 434 -1025 444 -1024
rect -43 -1068 35 -1026
rect -36 -1226 35 -1068
rect 95 -1226 105 -1026
rect 187 -1226 197 -1026
rect 252 -1226 262 -1026
rect 371 -1225 444 -1025
rect 496 -1225 506 -1024
rect 371 -1226 486 -1225
rect -36 -1227 79 -1226
<< via1 >>
rect 39 101 91 300
rect 195 100 251 301
rect 442 100 494 300
rect 276 10 328 62
rect 118 -162 170 -110
rect -49 -401 3 -200
rect 195 -400 251 -200
rect 356 -400 408 -199
rect -49 -728 3 -527
rect 195 -728 251 -528
rect 355 -728 407 -528
rect 117 -818 169 -766
rect 277 -985 329 -933
rect 35 -1226 95 -1026
rect 197 -1226 252 -1026
rect 444 -1225 496 -1024
<< metal2 >>
rect -44 345 494 386
rect -44 -190 -3 345
rect 35 301 95 311
rect 35 90 95 100
rect 195 301 251 311
rect 195 90 251 100
rect 442 300 494 345
rect 442 90 494 100
rect 276 62 328 72
rect 276 -24 328 10
rect 118 -76 328 -24
rect 118 -110 170 -76
rect 118 -172 170 -162
rect -49 -200 3 -190
rect -49 -411 3 -401
rect 195 -200 251 -190
rect 195 -410 251 -400
rect 355 -199 415 -189
rect 355 -410 415 -400
rect -44 -517 -3 -411
rect -49 -527 3 -517
rect -49 -738 3 -728
rect 195 -528 251 -518
rect 356 -519 416 -518
rect 195 -738 251 -728
rect 355 -528 416 -519
rect 355 -729 356 -728
rect 355 -737 416 -729
rect -44 -929 -3 -738
rect 356 -739 416 -737
rect 117 -766 169 -756
rect 117 -852 169 -818
rect 117 -904 329 -852
rect -46 -938 -3 -929
rect 277 -933 329 -904
rect -46 -995 -5 -938
rect 277 -995 329 -985
rect -44 -1004 -5 -995
rect -44 -1272 -3 -1004
rect 34 -1017 94 -1015
rect 34 -1025 95 -1017
rect 94 -1026 95 -1025
rect 27 -1226 34 -1216
rect 197 -1026 253 -1016
rect 95 -1226 103 -1216
rect 27 -1244 103 -1226
rect 197 -1236 253 -1226
rect 444 -1024 496 -1014
rect 444 -1235 496 -1225
rect 449 -1272 491 -1235
rect -44 -1313 491 -1272
<< via2 >>
rect 35 300 95 301
rect 35 101 39 300
rect 39 101 91 300
rect 91 101 95 300
rect 35 100 95 101
rect 195 100 251 301
rect 195 -400 251 -200
rect 355 -400 356 -199
rect 356 -400 408 -199
rect 408 -400 415 -199
rect 195 -728 251 -528
rect 356 -728 407 -528
rect 407 -728 416 -528
rect 356 -729 416 -728
rect 34 -1026 94 -1025
rect 34 -1226 35 -1026
rect 35 -1226 94 -1026
rect 197 -1226 252 -1026
rect 252 -1226 253 -1026
<< metal3 >>
rect 34 400 415 461
rect 34 306 95 400
rect 25 301 105 306
rect 25 100 35 301
rect 95 100 105 301
rect 25 95 105 100
rect 185 301 261 306
rect 185 100 195 301
rect 251 100 261 301
rect 185 95 261 100
rect 193 -195 253 95
rect 354 -194 415 400
rect 185 -200 261 -195
rect 185 -400 195 -200
rect 251 -400 261 -200
rect 185 -405 261 -400
rect 345 -199 425 -194
rect 345 -400 355 -199
rect 415 -400 425 -199
rect 345 -405 425 -400
rect 193 -523 253 -405
rect 354 -523 415 -405
rect 185 -528 261 -523
rect 185 -728 195 -528
rect 251 -728 261 -528
rect 185 -733 261 -728
rect 346 -528 426 -523
rect 346 -729 356 -528
rect 416 -729 426 -528
rect 32 -1020 93 -1019
rect 24 -1025 104 -1020
rect 194 -1021 255 -733
rect 346 -734 426 -729
rect 24 -1226 34 -1025
rect 94 -1226 104 -1025
rect 24 -1231 104 -1226
rect 187 -1026 263 -1021
rect 187 -1226 197 -1026
rect 253 -1226 263 -1026
rect 187 -1231 263 -1226
rect 32 -1326 93 -1231
rect 354 -1326 415 -734
rect 32 -1387 415 -1326
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729408613
transform 1 0 22 0 1 -1126
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729408613
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729408613
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729408613
transform 1 0 21 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729408613
transform 1 0 425 0 1 -300
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729408613
transform 1 0 21 0 1 -628
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729408613
transform 1 0 425 0 1 -628
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729408613
transform 1 0 426 0 1 -1126
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729408613
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729408613
transform 1 0 223 0 1 -300
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729408613
transform 1 0 223 0 1 -628
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729408613
transform 1 0 224 0 1 -1126
box -223 -200 223 200
<< labels >>
flabel viali 105 502 105 502 0 FreeSans 320 0 0 0 vdd
port 0 nsew
flabel metal3 65 425 65 425 0 FreeSans 320 0 0 0 d6
port 1 nsew
flabel metal1 142 -7 142 -7 0 FreeSans 320 0 0 0 vin
port 4 nsew
flabel metal1 426 234 426 234 0 FreeSans 320 0 0 0 out
port 8 nsew
flabel metal2 299 -917 299 -917 0 FreeSans 320 0 0 0 vpin
port 9 nsew
flabel metal3 224 -994 224 -994 0 FreeSans 320 0 0 0 d5
port 10 nsew
<< end >>
