magic
tech sky130A
magscale 1 2
timestamp 1729241942
<< psubdiff >>
rect -176 795 -106 829
rect 1042 795 1106 829
rect -176 756 -142 795
rect 1072 756 1106 795
rect -176 -110 -142 -67
rect 1072 -110 1106 -67
rect -176 -144 -106 -110
rect 1042 -144 1106 -110
<< psubdiffcont >>
rect -106 795 1042 829
rect -176 -67 -142 756
rect 1072 -67 1106 756
rect -106 -144 1042 -110
<< poly >>
rect -94 678 0 694
rect -94 644 -78 678
rect -44 644 0 678
rect -94 628 0 644
rect -30 623 0 628
rect 930 685 1022 701
rect 930 651 972 685
rect 1006 651 1022 685
rect 930 635 1022 651
rect 930 624 960 635
rect -30 56 0 88
rect -92 40 0 56
rect -92 6 -76 40
rect -42 6 0 40
rect -92 -10 0 6
rect 930 30 960 62
rect 930 14 1022 30
rect 930 -20 972 14
rect 1006 -20 1022 14
rect 930 -36 1022 -20
<< polycont >>
rect -78 644 -44 678
rect 972 651 1006 685
rect -76 6 -42 40
rect 972 -20 1006 14
<< locali >>
rect -176 795 -106 829
rect 1042 795 1106 829
rect -176 756 -142 795
rect 1072 756 1106 795
rect 972 685 1006 686
rect -94 644 -78 678
rect -44 644 -28 678
rect 956 651 972 685
rect 1006 651 1022 685
rect -79 627 -34 644
rect 962 634 1007 651
rect -76 567 -41 627
rect 969 624 1006 634
rect 972 568 1006 624
rect -76 67 -42 88
rect -76 57 -39 67
rect -77 40 -32 57
rect 972 41 1006 104
rect -92 6 -76 40
rect -42 6 -26 40
rect 969 31 1006 41
rect 962 14 1007 31
rect -76 5 -42 6
rect 956 -20 972 14
rect 1006 -20 1022 14
rect 972 -21 1006 -20
rect -176 -110 -142 -67
rect 275 -110 280 -109
rect 1072 -110 1106 -67
rect -176 -144 -106 -110
rect 1042 -144 1106 -110
<< viali >>
rect 220 829 272 838
rect 220 795 272 829
rect 658 795 717 829
rect 220 786 272 795
rect -78 644 -44 678
rect 972 651 1006 685
rect -76 6 -42 40
rect 972 -20 1006 14
rect 219 -110 275 -88
rect 657 -110 713 -99
rect 219 -144 275 -110
rect 657 -144 713 -110
rect 657 -155 713 -144
<< metal1 >>
rect 208 838 284 844
rect 208 786 220 838
rect 272 786 284 838
rect 646 829 661 835
rect 713 829 729 835
rect 646 795 658 829
rect 717 795 729 829
rect 646 789 661 795
rect 208 780 284 786
rect 651 783 661 789
rect 713 789 729 795
rect 713 783 723 789
rect 960 685 1018 691
rect -90 678 -32 684
rect -90 644 -78 678
rect -44 644 -30 678
rect 958 651 972 685
rect 1006 651 1018 685
rect 959 645 1018 651
rect -90 638 -31 644
rect -83 627 -31 638
rect 959 634 1011 645
rect -80 599 -38 627
rect -82 597 -36 599
rect -7 597 65 599
rect -82 399 65 597
rect 211 410 221 586
rect 273 410 283 586
rect -82 366 -36 399
rect -7 397 65 399
rect 429 397 439 599
rect 492 397 502 599
rect 969 598 1008 634
rect 647 398 657 598
rect 709 398 719 598
rect 865 399 1012 598
rect 865 398 937 399
rect 966 366 1012 399
rect -82 320 1012 366
rect -10 288 0 290
rect -73 88 0 288
rect 54 88 64 290
rect 211 88 221 289
rect 273 88 283 289
rect 442 88 488 320
rect 647 88 657 289
rect 709 88 719 289
rect 866 88 876 290
rect 928 289 938 290
rect 928 288 1002 289
rect 928 88 1012 288
rect -78 57 -39 88
rect -81 46 -29 57
rect -88 40 -29 46
rect -88 6 -76 40
rect -42 6 -28 40
rect 966 32 1012 88
rect 961 31 1012 32
rect 959 20 1012 31
rect 959 14 1018 20
rect -88 0 -30 6
rect 958 -20 972 14
rect 1006 -20 1018 14
rect 960 -26 1018 -20
rect 207 -88 287 -82
rect 207 -144 219 -88
rect 275 -144 287 -88
rect 207 -150 287 -144
rect 645 -99 725 -93
rect 645 -155 657 -99
rect 713 -155 725 -99
rect 645 -161 725 -155
<< via1 >>
rect 220 786 272 838
rect 661 829 713 835
rect 661 795 713 829
rect 661 783 713 795
rect 221 410 273 586
rect 439 397 492 599
rect 657 398 709 598
rect 0 88 54 290
rect 221 88 273 289
rect 657 88 709 289
rect 876 88 928 290
rect 219 -144 275 -88
rect 657 -155 713 -99
<< metal2 >>
rect 218 841 274 851
rect 218 775 274 785
rect 659 837 715 847
rect 659 771 715 781
rect 2 691 926 743
rect 2 397 54 691
rect 442 609 489 691
rect 219 598 275 608
rect 3 300 55 397
rect 219 387 275 397
rect 439 599 492 609
rect 439 387 492 397
rect 657 598 713 608
rect 657 388 713 398
rect 874 398 926 691
rect 0 291 55 300
rect 0 290 54 291
rect 0 4 54 88
rect 219 289 275 299
rect 219 78 275 88
rect 657 289 713 299
rect 874 291 928 398
rect 874 290 929 291
rect 657 78 713 88
rect 875 88 876 290
rect 928 88 929 290
rect 875 4 929 88
rect 0 -50 930 4
rect 219 -88 275 -78
rect 219 -162 275 -152
rect 657 -99 713 -89
rect 657 -165 713 -155
<< via2 >>
rect 218 838 274 841
rect 218 786 220 838
rect 220 786 272 838
rect 272 786 274 838
rect 218 785 274 786
rect 659 835 715 837
rect 659 783 661 835
rect 661 783 713 835
rect 713 783 715 835
rect 659 781 715 783
rect 219 586 275 598
rect 219 410 221 586
rect 221 410 273 586
rect 273 410 275 586
rect 219 397 275 410
rect 657 398 709 598
rect 709 398 713 598
rect 219 88 221 289
rect 221 88 273 289
rect 273 88 275 289
rect 657 88 709 289
rect 709 88 713 289
rect 219 -144 275 -96
rect 219 -152 275 -144
rect 657 -155 713 -99
<< metal3 >>
rect 208 841 284 846
rect 208 785 218 841
rect 274 785 284 841
rect 208 780 284 785
rect 649 837 725 842
rect 649 781 659 837
rect 715 781 725 837
rect 215 603 277 780
rect 649 776 725 781
rect 657 603 717 776
rect 209 598 285 603
rect 209 397 219 598
rect 275 397 285 598
rect 209 392 285 397
rect 647 598 723 603
rect 647 398 657 598
rect 713 398 723 598
rect 647 393 723 398
rect 209 289 285 294
rect 209 88 219 289
rect 275 88 285 289
rect 209 83 285 88
rect 647 289 723 294
rect 647 88 657 289
rect 713 88 723 289
rect 647 83 723 88
rect 216 -91 278 83
rect 209 -96 285 -91
rect 655 -94 716 83
rect 209 -152 219 -96
rect 275 -152 285 -96
rect 209 -157 285 -152
rect 647 -99 723 -94
rect 647 -155 657 -99
rect 713 -155 723 -99
rect 647 -160 723 -155
use sky130_fd_pr__nfet_01v8_6MBC9T  sky130_fd_pr__nfet_01v8_6MBC9T_0
timestamp 1729226061
transform 1 0 683 0 1 188
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_6MBC9T  sky130_fd_pr__nfet_01v8_6MBC9T_1
timestamp 1729226061
transform 1 0 247 0 1 188
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_6MBC9T  sky130_fd_pr__nfet_01v8_6MBC9T_2
timestamp 1729226061
transform 1 0 247 0 1 498
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_6MBC9T  sky130_fd_pr__nfet_01v8_6MBC9T_3
timestamp 1729226061
transform 1 0 683 0 1 498
box -247 -188 247 188
use sky130_fd_pr__nfet_01v8_SJFSNB  sky130_fd_pr__nfet_01v8_SJFSNB_0
timestamp 1729232893
transform 1 0 945 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_SJFSNB  sky130_fd_pr__nfet_01v8_SJFSNB_1
timestamp 1729232893
transform 1 0 -15 0 1 498
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_SJFSNB  sky130_fd_pr__nfet_01v8_SJFSNB_2
timestamp 1729232893
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_SJFSNB  sky130_fd_pr__nfet_01v8_SJFSNB_3
timestamp 1729232893
transform 1 0 945 0 1 498
box -73 -126 73 126
<< labels >>
flabel metal2 792 702 811 721 0 FreeSans 480 0 0 0 d9
port 0 nsew
flabel metal3 687 754 689 756 0 FreeSans 480 0 0 0 gnd
port 1 nsew
flabel metal1 980 340 982 342 0 FreeSans 480 0 0 0 d8
port 2 nsew
<< end >>
